----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06/07/2023 07:50:46 PM
-- Design Name: 
-- Module Name: Add_Subtract_4bit - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Add_Subtract_4bit is
    Port ( A0 : in STD_LOGIC;
           A1 : in STD_LOGIC;
           A2 : in STD_LOGIC;
           A3 : in STD_LOGIC;
           B0 : in STD_LOGIC;
           B1 : in STD_LOGIC;
           B2 : in STD_LOGIC;
           B3 : in STD_LOGIC;
           S0 : out STD_LOGIC;
           S1 : out STD_LOGIC;
           S2 : out STD_LOGIC;
           S3 : out STD_LOGIC;
           Overflow : out STD_LOGIC;
           Zero : out STD_LOGIC;
           CTR : in STD_LOGIC);
end Add_Subtract_4bit;
architecture Behavioral of Add_Subtract_4bit is
component FA
 port (
 A: in std_logic;
 B: in std_logic;
 C_in: in std_logic;
 S: out std_logic;
 C_out: out std_logic);
 end component;
 SIGNAL FA0_S, FA0_C, FA1_S, FA1_C, FA2_S, FA2_C, FA3_S, FA3_C, Bmod_0, Bmod_1, Bmod_2, Bmod_3  : std_logic;
 SIGNAL IS0 , IS1 , IS2 , IS3 : std_logic;
begin
 FA_0 : FA
 port map (
 A => A0,
 B => Bmod_0,
 C_in => CTR, -- Set to ground
 S => IS0,
 C_out => FA0_C);
 FA_1 : FA
 port map (
 A => A1,
 B => Bmod_1,
 C_in => FA0_C,
 S =>IS1,
 C_out => FA1_C);
 FA_2 : FA
 port map (
 A => A2,
 B => Bmod_2,
 C_in => FA1_C,
 S => IS2,
 C_out => FA2_C);
 FA_3 : FA
 port map (
 A => A3,
 B => Bmod_3,
 C_in => FA2_C,
 S => IS3,
 C_out => Overflow);
 
 Bmod_0 <= B0 XOR CTR;
 Bmod_1 <= B1 XOR CTR;
 Bmod_2 <= B2 XOR CTR;
 Bmod_3 <= B3 XOR CTR;
 S0 <= IS0;
 S1 <= IS1;
 S2 <= IS2;
 S3 <= IS3;
 Zero <= NOT(IS0 OR IS1 OR IS2 OR IS3);
end Behavioral;
----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06/07/2023 07:55:54 PM
-- Design Name: 
-- Module Name: Adder_3bit - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Adder_3bit is
    Port ( A0 : in STD_LOGIC;
           A1 : in STD_LOGIC;
           A2 : in STD_LOGIC;
           --B : in STD_LOGIC; -- Changed newly added
           S0 : out STD_LOGIC;
           S1 : out STD_LOGIC;
           S2 : out STD_LOGIC);
           --C_out : out STD_LOGIC);
           
           
end Adder_3bit;
architecture Behavioral of Adder_3bit is
component FA
 port (
 A: in std_logic;
 B: in std_logic :='0';
 C_in: in std_logic;
 S: out std_logic;
 C_out: out std_logic);
 end component;
 SIGNAL FA0_S, FA0_C, FA1_S, FA1_C, FA2_S, FA2_C, FA3_S, FA3_C  : std_logic;
begin
 FA_0 : FA
 port map (
 A => A0,
 --B => B, -- changed from 1 to 0
 C_in => '1', -- Set to ground
 S => S0,
 C_out => FA0_C);
 FA_1 : FA
 port map (
 A => A1,
 --B => '0',
 C_in => FA0_C,
 S => S1,
 C_out => FA1_C);
 FA_2 : FA
 port map (
 A => A2,
 --B => '0',
 C_in => FA1_C,
 S => S2);
 --C_out => FA2_C);
 
 

end Behavioral;